// Generator : SpinalHDL v1.4.2    git head : 804c7bd7b7feaddcc1d25ecef6c208fd5f776f79
// Component : cal_vn_serial
// Git hash  : f043fedd7462a55e48ae514eae5ce1768afb8b9c


module cal_vn_serial (
  input               en,
  input               vin_vld,
  input      [7:0]    v_in_0,
  input      [7:0]    v_in_1,
  input      [7:0]    v_in_2,
  input      [7:0]    v_in_3,
  input      [7:0]    v_in_4,
  input      [7:0]    v_in_5,
  input      [7:0]    v_in_6,
  input      [7:0]    v_in_7,
  output     [7:0]    vn_0,
  output     [7:0]    vn_1,
  output     [7:0]    vn_2,
  output     [7:0]    vn_3,
  output     [7:0]    vn_4,
  output     [7:0]    vn_5,
  output     [7:0]    vn_6,
  output     [7:0]    vn_7,
  output              vn_vld,
  input               clk,
  input               resetn
);
  wire       [11:0]   _zz_1;
  wire       [11:0]   _zz_2;
  wire       [11:0]   _zz_3;
  wire       [11:0]   _zz_4;
  wire       [11:0]   _zz_5;
  wire       [11:0]   _zz_6;
  wire       [11:0]   _zz_7;
  wire       [11:0]   _zz_8;
  reg        [7:0]    _zz_9;
  wire       [7:0]    FloorWrapVn_0_dout;
  wire       [7:0]    FloorWrapVn_1_dout;
  wire       [7:0]    FloorWrapVn_2_dout;
  wire       [7:0]    FloorWrapVn_3_dout;
  wire       [7:0]    FloorWrapVn_4_dout;
  wire       [7:0]    FloorWrapVn_5_dout;
  wire       [7:0]    FloorWrapVn_6_dout;
  wire       [7:0]    FloorWrapVn_7_dout;
  wire       [10:0]   _zz_10;
  wire       [11:0]   _zz_11;
  wire       [11:0]   _zz_12;
  wire       [11:0]   _zz_13;
  wire       [11:0]   _zz_14;
  wire       [11:0]   _zz_15;
  wire       [11:0]   _zz_16;
  wire       [11:0]   _zz_17;
  wire       [11:0]   _zz_18;
  wire       [11:0]   _zz_19;
  wire       [11:0]   _zz_20;
  wire       [11:0]   _zz_21;
  wire       [11:0]   _zz_22;
  wire       [11:0]   _zz_23;
  wire       [11:0]   _zz_24;
  wire       [11:0]   _zz_25;
  wire       [11:0]   _zz_26;
  reg                 in_vld_dly1;
  reg                 in_vld_dly2;
  reg        [2:0]    sum_cnt;
  reg                 sum_en;
  wire                sum_start;
  wire                sum_finish;
  reg        [10:0]   SumXinReg;
  wire       [10:0]   vin_ext_0;
  wire       [10:0]   vin_ext_1;
  wire       [10:0]   vin_ext_2;
  wire       [10:0]   vin_ext_3;
  wire       [10:0]   vin_ext_4;
  wire       [10:0]   vin_ext_5;
  wire       [10:0]   vin_ext_6;
  wire       [10:0]   vin_ext_7;
  wire       [11:0]   VinMinusMean_0;
  wire       [11:0]   VinMinusMean_1;
  wire       [11:0]   VinMinusMean_2;
  wire       [11:0]   VinMinusMean_3;
  wire       [11:0]   VinMinusMean_4;
  wire       [11:0]   VinMinusMean_5;
  wire       [11:0]   VinMinusMean_6;
  wire       [11:0]   VinMinusMean_7;
  wire       [7:0]    Vn_floor_0;
  wire       [7:0]    Vn_floor_1;
  wire       [7:0]    Vn_floor_2;
  wire       [7:0]    Vn_floor_3;
  wire       [7:0]    Vn_floor_4;
  wire       [7:0]    Vn_floor_5;
  wire       [7:0]    Vn_floor_6;
  wire       [7:0]    Vn_floor_7;
  reg        [7:0]    VnReg_0;
  reg        [7:0]    VnReg_1;
  reg        [7:0]    VnReg_2;
  reg        [7:0]    VnReg_3;
  reg        [7:0]    VnReg_4;
  reg        [7:0]    VnReg_5;
  reg        [7:0]    VnReg_6;
  reg        [7:0]    VnReg_7;

  assign _zz_10 = {{3{_zz_9[7]}}, _zz_9};
  assign _zz_11 = {vin_ext_0[10],vin_ext_0};
  assign _zz_12 = {SumXinReg[10],SumXinReg};
  assign _zz_13 = {vin_ext_1[10],vin_ext_1};
  assign _zz_14 = {SumXinReg[10],SumXinReg};
  assign _zz_15 = {vin_ext_2[10],vin_ext_2};
  assign _zz_16 = {SumXinReg[10],SumXinReg};
  assign _zz_17 = {vin_ext_3[10],vin_ext_3};
  assign _zz_18 = {SumXinReg[10],SumXinReg};
  assign _zz_19 = {vin_ext_4[10],vin_ext_4};
  assign _zz_20 = {SumXinReg[10],SumXinReg};
  assign _zz_21 = {vin_ext_5[10],vin_ext_5};
  assign _zz_22 = {SumXinReg[10],SumXinReg};
  assign _zz_23 = {vin_ext_6[10],vin_ext_6};
  assign _zz_24 = {SumXinReg[10],SumXinReg};
  assign _zz_25 = {vin_ext_7[10],vin_ext_7};
  assign _zz_26 = {SumXinReg[10],SumXinReg};
  FloorAndWrap FloorWrapVn_0 (
    .din     (_zz_1[11:0]              ), //i
    .dout    (FloorWrapVn_0_dout[7:0]  )  //o
  );
  FloorAndWrap FloorWrapVn_1 (
    .din     (_zz_2[11:0]              ), //i
    .dout    (FloorWrapVn_1_dout[7:0]  )  //o
  );
  FloorAndWrap FloorWrapVn_2 (
    .din     (_zz_3[11:0]              ), //i
    .dout    (FloorWrapVn_2_dout[7:0]  )  //o
  );
  FloorAndWrap FloorWrapVn_3 (
    .din     (_zz_4[11:0]              ), //i
    .dout    (FloorWrapVn_3_dout[7:0]  )  //o
  );
  FloorAndWrap FloorWrapVn_4 (
    .din     (_zz_5[11:0]              ), //i
    .dout    (FloorWrapVn_4_dout[7:0]  )  //o
  );
  FloorAndWrap FloorWrapVn_5 (
    .din     (_zz_6[11:0]              ), //i
    .dout    (FloorWrapVn_5_dout[7:0]  )  //o
  );
  FloorAndWrap FloorWrapVn_6 (
    .din     (_zz_7[11:0]              ), //i
    .dout    (FloorWrapVn_6_dout[7:0]  )  //o
  );
  FloorAndWrap FloorWrapVn_7 (
    .din     (_zz_8[11:0]              ), //i
    .dout    (FloorWrapVn_7_dout[7:0]  )  //o
  );
  always @(*) begin
    case(sum_cnt)
      3'b000 : begin
        _zz_9 = v_in_0;
      end
      3'b001 : begin
        _zz_9 = v_in_1;
      end
      3'b010 : begin
        _zz_9 = v_in_2;
      end
      3'b011 : begin
        _zz_9 = v_in_3;
      end
      3'b100 : begin
        _zz_9 = v_in_4;
      end
      3'b101 : begin
        _zz_9 = v_in_5;
      end
      3'b110 : begin
        _zz_9 = v_in_6;
      end
      default : begin
        _zz_9 = v_in_7;
      end
    endcase
  end

  assign sum_start = (sum_cnt == 3'b000);
  assign sum_finish = (sum_cnt == 3'b111);
  assign vin_ext_0 = {v_in_0,3'b000};
  assign vin_ext_1 = {v_in_1,3'b000};
  assign vin_ext_2 = {v_in_2,3'b000};
  assign vin_ext_3 = {v_in_3,3'b000};
  assign vin_ext_4 = {v_in_4,3'b000};
  assign vin_ext_5 = {v_in_5,3'b000};
  assign vin_ext_6 = {v_in_6,3'b000};
  assign vin_ext_7 = {v_in_7,3'b000};
  assign VinMinusMean_0 = ($signed(_zz_11) - $signed(_zz_12));
  assign VinMinusMean_1 = ($signed(_zz_13) - $signed(_zz_14));
  assign VinMinusMean_2 = ($signed(_zz_15) - $signed(_zz_16));
  assign VinMinusMean_3 = ($signed(_zz_17) - $signed(_zz_18));
  assign VinMinusMean_4 = ($signed(_zz_19) - $signed(_zz_20));
  assign VinMinusMean_5 = ($signed(_zz_21) - $signed(_zz_22));
  assign VinMinusMean_6 = ($signed(_zz_23) - $signed(_zz_24));
  assign VinMinusMean_7 = ($signed(_zz_25) - $signed(_zz_26));
  assign _zz_1 = VinMinusMean_0;
  assign Vn_floor_0 = FloorWrapVn_0_dout;
  assign _zz_2 = VinMinusMean_1;
  assign Vn_floor_1 = FloorWrapVn_1_dout;
  assign _zz_3 = VinMinusMean_2;
  assign Vn_floor_2 = FloorWrapVn_2_dout;
  assign _zz_4 = VinMinusMean_3;
  assign Vn_floor_3 = FloorWrapVn_3_dout;
  assign _zz_5 = VinMinusMean_4;
  assign Vn_floor_4 = FloorWrapVn_4_dout;
  assign _zz_6 = VinMinusMean_5;
  assign Vn_floor_5 = FloorWrapVn_5_dout;
  assign _zz_7 = VinMinusMean_6;
  assign Vn_floor_6 = FloorWrapVn_6_dout;
  assign _zz_8 = VinMinusMean_7;
  assign Vn_floor_7 = FloorWrapVn_7_dout;
  assign vn_0 = VnReg_0;
  assign vn_1 = VnReg_1;
  assign vn_2 = VnReg_2;
  assign vn_3 = VnReg_3;
  assign vn_4 = VnReg_4;
  assign vn_5 = VnReg_5;
  assign vn_6 = VnReg_6;
  assign vn_7 = VnReg_7;
  assign vn_vld = (sum_finish && sum_en);
  always @ (posedge clk or negedge resetn) begin
    if (!resetn) begin
      in_vld_dly1 <= 1'b0;
      in_vld_dly2 <= 1'b0;
      sum_cnt <= 3'b000;
      sum_en <= 1'b0;
      SumXinReg <= 11'h0;
      VnReg_0 <= 8'h0;
      VnReg_1 <= 8'h0;
      VnReg_2 <= 8'h0;
      VnReg_3 <= 8'h0;
      VnReg_4 <= 8'h0;
      VnReg_5 <= 8'h0;
      VnReg_6 <= 8'h0;
      VnReg_7 <= 8'h0;
    end else begin
      if(en)begin
        in_vld_dly1 <= vin_vld;
        in_vld_dly2 <= in_vld_dly1;
      end else begin
        in_vld_dly1 <= 1'b0;
        in_vld_dly2 <= 1'b0;
      end
      if(en)begin
        if(vin_vld)begin
          sum_en <= 1'b1;
        end else begin
          if(sum_finish)begin
            sum_en <= 1'b0;
          end
        end
      end else begin
        sum_en <= 1'b0;
      end
      if(sum_en)begin
        sum_cnt <= (sum_cnt + 3'b001);
        if(sum_start)begin
          SumXinReg <= {{3{v_in_0[7]}}, v_in_0};
        end else begin
          SumXinReg <= ($signed(SumXinReg) + $signed(_zz_10));
        end
      end else begin
        sum_cnt <= 3'b000;
      end
      if((sum_finish && sum_en))begin
        VnReg_0 <= Vn_floor_0;
        VnReg_1 <= Vn_floor_1;
        VnReg_2 <= Vn_floor_2;
        VnReg_3 <= Vn_floor_3;
        VnReg_4 <= Vn_floor_4;
        VnReg_5 <= Vn_floor_5;
        VnReg_6 <= Vn_floor_6;
        VnReg_7 <= Vn_floor_7;
      end
    end
  end


endmodule
